/*
*   Copyright 2016 Purdue University
*
*   Licensed under the Apache License, Version 2.0 (the "License");
*   you may not use this file except in compliance with the License.
*   You may obtain a copy of the License at
*
*       http://www.apache.org/licenses/LICENSE-2.0
*
*   Unless required by applicable law or agreed to in writing, software
*   distributed under the License is distributed on an "AS IS" BASIS,
*   WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
*   See the License for the specific language governing permissions and
*   limitations under the License.
*
*
*   Filename:     cpu_tracker.sv
*
*   Created by:   Jacob R. Stevens
*   Email:        steven69@purdue.edu
*   Date Created: 06/27/2016
*   Description:  Prints out a trace of the cpu executing that can be
*                 compared against the trace generated by the ISS

    Updated by:   Anusyua Nallathambi, Ansh Patel, Zach Lagpacan
    Date: 10/21/2024
*/

`include "cpu_types_pkg.vh"
import cpu_types_pkg::*;

module cpu_tracker_rv32(
  input logic CLK,
  input logic wb_stall,
  input logic dhit,
  input logic[FUNC3_W-1:0] funct_3,
  input logic[FUNC7_W-1:0] funct_7,
  input opcode_t opcode,
  input regbits_t rs1,
  input regbits_t rs2,
  input regbits_t wsel,
  input word_t instr,
  input word_t pc,
  input word_t next_pc_val,
  input word_t branch_addr,
  input word_t jump_addr,
  input word_t imm,
  input logic [19:0] lui_pre_shift,
  input word_t store_dat,
  input word_t reg_dat,
  input word_t load_dat,
  input word_t dat_addr
);

  parameter CPUID = 1;

  integer fptr, halt_written;
  string filename;
  string instr_mnemonic, output_str, operands, temp_str, halt_temp_str;
  string rs1_str, rs2_str, ram_str, lw_str, halt_output_str, dest_str;
  opcode_t last_opcode;
  funct3_r_t funct3_r;
  funct3_i_t funct3_i;
  funct3_ld_i_t funct3_ld_i;
  funct3_s_t funct3_s;
  funct7_r_t funct7_r;
  funct7_srla_r_t funct7_srla_r;
  funct3_b_t funct3_b;

  string upper_instr;
  string upper_pc;
  string upper_next_pc_val;
  string upper_lui;
  string upper_auipc;
  string upper_store_dat;
  string upper_reg_dat;
  string upper_load_dat;
  string upper_dat_addr;

  word_t presumed_reserve_addr;
  string upper_presumed_reserve_addr;

  initial begin: INIT_FILE
    $sformat(filename, "cpu%0d_trace.log", CPUID);
		fptr = $fopen(filename, "w");
    halt_written = 0;
  end

  always_comb begin
    rs1_str    = registerAssign(rs1);
    rs2_str    = registerAssign(rs2);
    dest_str  = registerAssign(wsel);
  end

  always_comb begin
    case (opcode)
      RTYPE: $sformat(operands, "%s, %s, %s", dest_str, rs1_str, rs2_str);
      ITYPE: 
      begin
        case(funct3_i_t'(funct_3))
          SRLI_SRAI, SLLI: $sformat(operands, "%s, %s, %0d", dest_str, rs1_str, (imm[4:0]));
          default: $sformat(operands, "%s, %s, %0d", dest_str, rs1_str, signed'(imm));
        endcase
      end
      ITYPE_LW: $sformat(operands, "%s, %0d(%s)", dest_str, signed'(imm), rs1_str);
      LR_SC:
      begin
        case(funct5_atomic_t'(funct_7[6:2]))
          LR: $sformat(operands, "%s, (%s)", dest_str, rs1_str);
          SC: $sformat(operands, "%s, %s, (%s)", dest_str, rs2_str, rs1_str);
        endcase
      end
      STYPE: $sformat(operands, "%s, %0d(%s)", rs2_str, signed'(imm), rs1_str);
      JALR: $sformat(operands, "%s, %s, %0d", dest_str, rs1_str, signed'(imm));
      BTYPE: $sformat(operands, "%s, %s, %0d", rs1_str, rs2_str, signed'(branch_addr));
      JAL: $sformat(operands, "%s, %0d", dest_str, signed'(jump_addr));
      LUI:   $sformat(operands,"%s, %0d", dest_str, signed'(lui_pre_shift));
      AUIPC: $sformat(operands,"%s, %0d", dest_str, signed'(lui_pre_shift));
      HALT:  $sformat(operands, "");
    endcase
  end

  always_comb begin
    case (opcode)
      JAL:      instr_mnemonic = "JAL";
      JALR:      instr_mnemonic = "JALR";
      BTYPE:
      begin
        case(funct3_b_t'(funct_3))
          BEQ:      instr_mnemonic = "BEQ";
          BNE:      instr_mnemonic = "BNE";
          BLT:      instr_mnemonic = "BLT";
          BGE:      instr_mnemonic = "BGE";
          BLTU:     instr_mnemonic = "BLTU";
          BGEU:     instr_mnemonic = "BGEU";
        endcase
      end
      STYPE:
      begin
        case(funct3_s_t'(funct_3))
          SB:       instr_mnemonic = "SB";
          SH:       instr_mnemonic = "SH";
          SW:       instr_mnemonic = "SW";
        endcase
      end
      ITYPE_LW:
      begin
        case(funct3_ld_i_t'(funct_3))
          LB:       instr_mnemonic = "LB";
          LH:       instr_mnemonic = "LH";
          LW:       instr_mnemonic = "LW";
          LBU:      instr_mnemonic = "LBU";
          LHU:      instr_mnemonic = "LHU";
        endcase
      end
      LR_SC:
      begin
        case(funct5_atomic_t'(funct_7[6:2]))
          LR:       instr_mnemonic = "LR.W";
          SC:       instr_mnemonic = "SC.W";
        endcase
      end
      ITYPE:
      begin
        case(funct3_i_t'(funct_3))
          ADDI:     instr_mnemonic = "ADDI";
          SLTI:     instr_mnemonic = "SLTI";
          SLTIU:    instr_mnemonic = "SLTIU";
          ANDI:     instr_mnemonic = "ANDI";
          ORI:      instr_mnemonic = "ORI";
          XORI:     instr_mnemonic = "XORI";
          SLLI:     instr_mnemonic = "SLLI";
          SRLI_SRAI:    
          begin
            case(funct7_srla_r_t'(funct_7))
              SRA: instr_mnemonic = "SRAI";
              SRL: instr_mnemonic = "SRLI";
            endcase
          end
        endcase
      end
      LUI:      instr_mnemonic = "LUI";
      AUIPC:   instr_mnemonic = "AUIPC";
      HALT:     instr_mnemonic = "HALT";
      RTYPE: begin
        case(funct3_r_t'(funct_3))
          SLL:  instr_mnemonic = "SLL";
          SRL_SRA:
          begin
            case(funct7_srla_r_t'(funct_7))
              SRA: instr_mnemonic = "SRA";
              SRL: instr_mnemonic = "SRL";
            endcase
          end
          ADD_SUB:  
          begin
            case(funct7_r_t'(funct_7))
              ADD: instr_mnemonic = "ADD";
              SUB: instr_mnemonic = "SUB";
            endcase
          end
          AND:  instr_mnemonic = "AND";
          OR:   instr_mnemonic = "OR";
          XOR:  instr_mnemonic = "XOR";
          SLT:  instr_mnemonic = "SLT";
          SLTU: instr_mnemonic = "SLTU";
        endcase
      end
      default:  instr_mnemonic = "xxx";
    endcase
  end

  function string registerAssign(input logic [4:0] register);
    case (register)
      5'd0:   registerAssign = "R0";
      5'd1:   registerAssign = "R1";
      5'd2:   registerAssign = "R2";
      5'd3:   registerAssign = "R3";
      5'd4:   registerAssign = "R4";
      5'd5:   registerAssign = "R5";
      5'd6:   registerAssign = "R6";
      5'd7:   registerAssign = "R7";
      5'd8:   registerAssign = "R8";
      5'd9:   registerAssign = "R9";
      5'd10:  registerAssign = "R10";
      5'd11:  registerAssign = "R11";
      5'd12:  registerAssign = "R12";
      5'd13:  registerAssign = "R13";
      5'd14:  registerAssign = "R14";
      5'd15:  registerAssign = "R15";
      5'd16:  registerAssign = "R16";
      5'd17:  registerAssign = "R17";
      5'd18:  registerAssign = "R18";
      5'd19:  registerAssign = "R19";
      5'd20:  registerAssign = "R20";
      5'd21:  registerAssign = "R21";
      5'd22:  registerAssign = "R22";
      5'd23:  registerAssign = "R23";
      5'd24:  registerAssign = "R24";
      5'd25:  registerAssign = "R25";
      5'd26:  registerAssign = "R26";
      5'd27:  registerAssign = "R27";
      5'd28:  registerAssign = "R28";
      5'd29:  registerAssign = "R29";
      5'd30:  registerAssign = "R30";
      5'd31:  registerAssign = "R31";
    endcase
  endfunction

  // always_ff @ (posedge CLK) begin
    // if (dhit) begin
        // if (last_opcode == ITYPE_LW) begin
        // if (opcode == ITYPE_LW) begin
        //   $sformat(temp_str, "%X (Core %d): %X", pc, CPUID + 1, instr);
        //   $sformat(temp_str, "%s %s %s\n", temp_str, instr_mnemonic, operands);
        //   $sformat(ram_str, "    [word read");
        //   $sformat(ram_str, "%s from %x]\n", ram_str, {16'h0, dat_addr[15:0]});
        //   $sformat(ram_str, "%s    %s", ram_str, dest_str);
        //   $sformat(ram_str, "%s <-- %x\n", ram_str, load_dat);
        //   $sformat(lw_str, "%s%s\n", temp_str, ram_str);
        //   $fwrite(fptr, lw_str);
        // end
    // end
  // end

  always_ff @ (posedge CLK) begin
    if (!wb_stall)
      last_opcode <= opcode;
  end

  always_comb begin
    upper_instr = $sformatf("%X", instr);
    upper_instr = upper_instr.toupper();
    upper_pc = $sformatf("%X", pc);
    upper_pc = upper_pc.toupper();
    upper_next_pc_val = $sformatf("%X", next_pc_val);
    upper_next_pc_val = upper_next_pc_val.toupper();
    upper_lui = $sformatf("%X", {lui_pre_shift, 12'b0});
    upper_lui = upper_lui.toupper();
    upper_auipc = $sformatf("%X", pc+(lui_pre_shift<<12));
    upper_auipc = upper_auipc.toupper();
    upper_store_dat = $sformatf("%X", store_dat);
    upper_store_dat = upper_store_dat.toupper();
    upper_reg_dat = $sformatf("%X", reg_dat);
    upper_reg_dat = upper_reg_dat.toupper();
    upper_load_dat = $sformatf("%X", load_dat);
    upper_load_dat = upper_load_dat.toupper();
    upper_dat_addr = $sformatf("%X", {16'h0, dat_addr[15:0]});
    upper_dat_addr = upper_dat_addr.toupper();
    upper_presumed_reserve_addr = $sformatf("%X", presumed_reserve_addr + 32'h1);
    upper_presumed_reserve_addr = upper_presumed_reserve_addr.toupper();
  end

  always_ff @ (posedge CLK) begin
    if (!wb_stall && instr != 0 && instr != 32'h00000013) begin
      $sformat(temp_str, "%s(Core %0d): %s", upper_pc, CPUID, upper_instr);
      $sformat(temp_str, "%s %s %s\n", temp_str, instr_mnemonic, operands);
      $sformat(temp_str, "%s\tPC <-- %s\n", temp_str, upper_next_pc_val);
      case(opcode)
        RTYPE: 
        begin
          $sformat(temp_str, "%s\t%s <-- %s\n", temp_str, dest_str, upper_reg_dat);
        end
        ITYPE:
        begin
          case(funct3_i_t'(funct_3))
            default: $sformat(temp_str, "%s\t%s <-- %s\n", temp_str, dest_str, upper_reg_dat);
          endcase
        end
        BTYPE:
        begin
          // pass
        end
        JAL, JALR: $sformat(temp_str, "%s\t%s <-- %s\n", temp_str, dest_str, upper_reg_dat);
        LUI:  $sformat(temp_str, "%s\t%s <-- %s\n", temp_str, dest_str, upper_lui);
        AUIPC:  $sformat(temp_str, "%s\t%s <-- %s\n", temp_str, dest_str, upper_auipc);
        STYPE: begin
              $sformat(temp_str,"%s\t[%s]",temp_str,upper_dat_addr);
              $sformat(temp_str, "%s <-- %s\n", temp_str, upper_store_dat);
        end
        ITYPE_LW:
        begin
          $sformat(ram_str, "\t[word read");
          $sformat(ram_str, "%s from %s]\n", ram_str, upper_dat_addr);
          $sformat(ram_str, "%s\t%s", ram_str, dest_str);
          $sformat(ram_str, "%s <-- %s\n", ram_str, upper_load_dat);
          $sformat(temp_str, "%s%s", temp_str, ram_str);
        end
        LR_SC:
        begin
          case(funct5_atomic_t'(funct_7[6:2]))
            LR: begin
              $sformat(ram_str, "\t[word read");
              $sformat(ram_str, "%s from %s]\n", ram_str, upper_dat_addr);
              $sformat(ram_str, "%s\t%s", ram_str, dest_str);
              $sformat(ram_str, "%s <-- %s\n", ram_str, upper_load_dat);
              presumed_reserve_addr <= {dat_addr[31:1], 1'b0};
              $sformat(ram_str, "%s\tRMW <-- %s\n", ram_str, upper_dat_addr);
              $sformat(temp_str, "%s%s", temp_str, ram_str);
            end
            SC: begin
              if (reg_dat == 0) begin
                $sformat(temp_str,"%s\t[%s]",temp_str,upper_dat_addr);
                $sformat(temp_str, "%s <-- %s\n", temp_str, upper_store_dat);
              end
              $sformat(temp_str, "%s\t%s <-- %s\n", temp_str, dest_str, upper_reg_dat);
              if (reg_dat == 0) begin
                $sformat(temp_str, "%s\tRMW <-- %s\n", temp_str, upper_presumed_reserve_addr);
              end
            end
          endcase
        end
        default: $sformat(temp_str, "");
      endcase
      $sformat(output_str, "%s\n", temp_str);
      $fwrite(fptr, output_str);
    end
  end

  final begin: CLOSE_FILE
    $fclose(fptr);
  end

endmodule